module sort1(
  // Input signals
  N0, N1, N2, N3, N4, N5,
  // Output signals
  S0, S1, S2, S3, S4, S5 
);

input [5:0] N0, N1, N2, N3, N4, N5;

output reg S0, S1, S2, S3, S4, S5;

always @(*) begin
  if () begin
    
  end
  
end


endmodule