`timescale 1ns/100ps

module dummyModule();
endmodule


