 always @(posedge clk) begin

     b = a;

     c = b; //b,c同時
     
 end